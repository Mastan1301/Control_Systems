OPMODEL1.CIR - OPAMP MODEL SINGLE-POLE
*
VS	8	0	AC	1  SIN(0VOFF 1VPEAK   1KHZ)
XOP	1 0	3	OPAMP1
RS	8	1	100
RL	3	0	3.33K

* FEEDBACK LOOP
R2	3	7	9K
R1	7	0	1K

*
* OPAMP MACRO MODEL, SINGLE-POLE
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   output
*                   |   |   |
.SUBCKT OPAMP1	    1   2   6
* INPUT IMPEDANCE
RIN	1	7	1K
* DC GAIN=10K AND POLE AT 200KHz
EGAIN	3 0	1 2	10K
RP1	3	4	1K
CP1	4	0	31UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER	5 0	4 0	1
ROUT	5	6	10K
.ENDS
*
* ANALYSIS
.TRAN 	1US  100MS
*.PLOT	AC 	VM(3)
.PROBE
.END
